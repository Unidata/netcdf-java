netcdf writeEnumType {
  types:
    short enum dessertType { 'pie' = 18, 'donut' = 268, 'cake' = 3284};
    enum dessert { 'pie' = 18, 'donut' = 268, 'cake' = 3284};

  dimensions:
    time = UNLIMITED;   // (3 currently)
  variables:
    enum dessert dessert(time=3);
      :_ChunkSizes = 4096U; // uint

  // global attributes:

  data:
    dessert =
      {18, 268, 3284}
}